// Global nets module 

`celldefine
module cds_globals;


supply0 vss_;

supply1 vdd_;


endmodule
`endcelldefine
